library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity hex is
port (
    clk: in  std_logic;
    addr: in  std_logic_vector(15 downto 0);
    dout: out std_logic_vector(39 downto 0) := (others => '0')
    );
end hex;

architecture Behavioral of hex is
type CODE_ARRAY is array (NATURAL RANGE <>) OF std_logic_vector(39 downto 0);

constant MAX_CNT: integer := 651;
signal mem: CODE_ARRAY(MAX_CNT downto 0); 


begin
    
process(clk)
begin
if (clk' event and clk = '1') then
    dout <= mem(conv_integer(addr));
end if;
end process;


mem(0)<=x"2300000000";
mem(1)<=x"0200000012";
mem(2)<=x"2300070003";
mem(3)<=x"0200000012";
mem(4)<=x"2300000064";
mem(5)<=x"0200000024";
mem(6)<=x"23000003e8";
mem(7)<=x"0200000025";
mem(8)<=x"230000000a";
mem(9)<=x"0200000026";
mem(10)<=x"51000001c2";
mem(11)<=x"510000025e";
mem(12)<=x"2200000000";
mem(13)<=x"510000025e";
mem(14)<=x"2200000001";
mem(15)<=x"510000025e";
mem(16)<=x"2200000002";
mem(17)<=x"2100000001";
mem(18)<=x"3700000000";
mem(19)<=x"3700000000";
mem(20)<=x"3100000002";
mem(21)<=x"2200000003";
mem(22)<=x"0200000020";
mem(23)<=x"4100000020";
mem(24)<=x"0100000022";
mem(25)<=x"2200000004";
mem(26)<=x"2300000001";
mem(27)<=x"2200000005";
mem(28)<=x"2100000000";
mem(29)<=x"3400000005";
mem(30)<=x"1200000043";
mem(31)<=x"2300000002";
mem(32)<=x"2200000005";
mem(33)<=x"2100000000";
mem(34)<=x"3400000005";
mem(35)<=x"1200000045";
mem(36)<=x"2300000003";
mem(37)<=x"2200000005";
mem(38)<=x"2100000000";
mem(39)<=x"3400000005";
mem(40)<=x"1200000047";
mem(41)<=x"2300000011";
mem(42)<=x"2200000005";
mem(43)<=x"2100000000";
mem(44)<=x"3400000005";
mem(45)<=x"1200000049";
mem(46)<=x"2300000022";
mem(47)<=x"2200000005";
mem(48)<=x"2100000000";
mem(49)<=x"3400000005";
mem(50)<=x"120000004b";
mem(51)<=x"2300000050";
mem(52)<=x"2200000005";
mem(53)<=x"2100000000";
mem(54)<=x"3400000005";
mem(55)<=x"120000004d";
mem(56)<=x"2300000004";
mem(57)<=x"2200000005";
mem(58)<=x"2100000000";
mem(59)<=x"3400000005";
mem(60)<=x"120000004f";
mem(61)<=x"2300000099";
mem(62)<=x"2200000005";
mem(63)<=x"2100000000";
mem(64)<=x"3400000005";
mem(65)<=x"1200000051";
mem(66)<=x"1100000053";
mem(67)<=x"5100000055";
mem(68)<=x"110000000a";
mem(69)<=x"5100000059";
mem(70)<=x"110000000a";
mem(71)<=x"510000005d";
mem(72)<=x"110000000a";
mem(73)<=x"5100000061";
mem(74)<=x"110000000a";
mem(75)<=x"510000009c";
mem(76)<=x"110000000a";
mem(77)<=x"51000000d7";
mem(78)<=x"110000000a";
mem(79)<=x"5100000126";
mem(80)<=x"110000000a";
mem(81)<=x"510000019d";
mem(82)<=x"110000000a";
mem(83)<=x"5100000231";
mem(84)<=x"110000000a";
mem(85)<=x"2100000004";
mem(86)<=x"0200000024";
mem(87)<=x"5100000204";
mem(88)<=x"5200000000";
mem(89)<=x"2100000004";
mem(90)<=x"0200000025";
mem(91)<=x"5100000204";
mem(92)<=x"5200000000";
mem(93)<=x"2100000004";
mem(94)<=x"0200000026";
mem(95)<=x"5100000204";
mem(96)<=x"5200000000";
mem(97)<=x"2100000004";
mem(98)<=x"0200000027";
mem(99)<=x"2300000001";
mem(100)<=x"0200000028";
mem(101)<=x"4100000100";
mem(102)<=x"2300000000";
mem(103)<=x"0200000028";
mem(104)<=x"230000004f";
mem(105)<=x"0200000010";
mem(106)<=x"230000006e";
mem(107)<=x"0200000010";
mem(108)<=x"2300000065";
mem(109)<=x"0200000010";
mem(110)<=x"2300000050";
mem(111)<=x"0200000010";
mem(112)<=x"2300000075";
mem(113)<=x"0200000010";
mem(114)<=x"230000006c";
mem(115)<=x"0200000010";
mem(116)<=x"2300000073";
mem(117)<=x"0200000010";
mem(118)<=x"2300000065";
mem(119)<=x"0200000010";
mem(120)<=x"2300000020";
mem(121)<=x"0200000010";
mem(122)<=x"2300000054";
mem(123)<=x"0200000010";
mem(124)<=x"2300000065";
mem(125)<=x"0200000010";
mem(126)<=x"2300000073";
mem(127)<=x"0200000010";
mem(128)<=x"2300000074";
mem(129)<=x"0200000010";
mem(130)<=x"230000002e";
mem(131)<=x"0200000010";
mem(132)<=x"2300000020";
mem(133)<=x"0200000010";
mem(134)<=x"2300000050";
mem(135)<=x"0200000010";
mem(136)<=x"2300000077";
mem(137)<=x"0200000010";
mem(138)<=x"230000006d";
mem(139)<=x"0200000010";
mem(140)<=x"2300000020";
mem(141)<=x"0200000010";
mem(142)<=x"230000004e";
mem(143)<=x"0200000010";
mem(144)<=x"2300000075";
mem(145)<=x"0200000010";
mem(146)<=x"230000006d";
mem(147)<=x"0200000010";
mem(148)<=x"230000003a";
mem(149)<=x"0200000010";
mem(150)<=x"0100000027";
mem(151)<=x"5100000265";
mem(152)<=x"230000000a";
mem(153)<=x"0200000010";
mem(154)<=x"5100000204";
mem(155)<=x"5200000000";
mem(156)<=x"2100000004";
mem(157)<=x"0200000027";
mem(158)<=x"2300000002";
mem(159)<=x"0200000028";
mem(160)<=x"4100000100";
mem(161)<=x"2300000000";
mem(162)<=x"0200000028";
mem(163)<=x"2300000054";
mem(164)<=x"0200000010";
mem(165)<=x"2300000077";
mem(166)<=x"0200000010";
mem(167)<=x"230000006f";
mem(168)<=x"0200000010";
mem(169)<=x"2300000050";
mem(170)<=x"0200000010";
mem(171)<=x"2300000075";
mem(172)<=x"0200000010";
mem(173)<=x"230000006c";
mem(174)<=x"0200000010";
mem(175)<=x"2300000073";
mem(176)<=x"0200000010";
mem(177)<=x"2300000065";
mem(178)<=x"0200000010";
mem(179)<=x"2300000020";
mem(180)<=x"0200000010";
mem(181)<=x"2300000054";
mem(182)<=x"0200000010";
mem(183)<=x"2300000065";
mem(184)<=x"0200000010";
mem(185)<=x"2300000073";
mem(186)<=x"0200000010";
mem(187)<=x"2300000074";
mem(188)<=x"0200000010";
mem(189)<=x"230000002e";
mem(190)<=x"0200000010";
mem(191)<=x"2300000020";
mem(192)<=x"0200000010";
mem(193)<=x"2300000050";
mem(194)<=x"0200000010";
mem(195)<=x"2300000077";
mem(196)<=x"0200000010";
mem(197)<=x"230000006d";
mem(198)<=x"0200000010";
mem(199)<=x"2300000020";
mem(200)<=x"0200000010";
mem(201)<=x"230000004e";
mem(202)<=x"0200000010";
mem(203)<=x"2300000075";
mem(204)<=x"0200000010";
mem(205)<=x"230000006d";
mem(206)<=x"0200000010";
mem(207)<=x"230000003a";
mem(208)<=x"0200000010";
mem(209)<=x"0100000027";
mem(210)<=x"5100000265";
mem(211)<=x"230000000a";
mem(212)<=x"0200000010";
mem(213)<=x"5100000204";
mem(214)<=x"5200000000";
mem(215)<=x"2300000056";
mem(216)<=x"0200000010";
mem(217)<=x"2300000043";
mem(218)<=x"0200000010";
mem(219)<=x"2300000050";
mem(220)<=x"0200000010";
mem(221)<=x"2300000031";
mem(222)<=x"0200000010";
mem(223)<=x"230000003a";
mem(224)<=x"0200000010";
mem(225)<=x"010000002d";
mem(226)<=x"5100000265";
mem(227)<=x"230000000a";
mem(228)<=x"0200000010";
mem(229)<=x"2300000056";
mem(230)<=x"0200000010";
mem(231)<=x"2300000043";
mem(232)<=x"0200000010";
mem(233)<=x"2300000050";
mem(234)<=x"0200000010";
mem(235)<=x"2300000032";
mem(236)<=x"0200000010";
mem(237)<=x"230000003a";
mem(238)<=x"0200000010";
mem(239)<=x"010000002d";
mem(240)<=x"3800000000";
mem(241)<=x"3800000000";
mem(242)<=x"3800000000";
mem(243)<=x"3800000000";
mem(244)<=x"5100000265";
mem(245)<=x"230000000a";
mem(246)<=x"0200000010";
mem(247)<=x"2300000049";
mem(248)<=x"0200000010";
mem(249)<=x"2300000041";
mem(250)<=x"0200000010";
mem(251)<=x"2300000043";
mem(252)<=x"0200000010";
mem(253)<=x"2300000031";
mem(254)<=x"0200000010";
mem(255)<=x"230000003a";
mem(256)<=x"0200000010";
mem(257)<=x"010000002e";
mem(258)<=x"5100000265";
mem(259)<=x"230000000a";
mem(260)<=x"0200000010";
mem(261)<=x"2300000049";
mem(262)<=x"0200000010";
mem(263)<=x"2300000041";
mem(264)<=x"0200000010";
mem(265)<=x"2300000043";
mem(266)<=x"0200000010";
mem(267)<=x"2300000032";
mem(268)<=x"0200000010";
mem(269)<=x"230000003a";
mem(270)<=x"0200000010";
mem(271)<=x"010000002e";
mem(272)<=x"3800000000";
mem(273)<=x"3800000000";
mem(274)<=x"3800000000";
mem(275)<=x"3800000000";
mem(276)<=x"5100000265";
mem(277)<=x"230000000a";
mem(278)<=x"0200000010";
mem(279)<=x"2300000049";
mem(280)<=x"0200000010";
mem(281)<=x"2300000041";
mem(282)<=x"0200000010";
mem(283)<=x"2300000043";
mem(284)<=x"0200000010";
mem(285)<=x"2300000033";
mem(286)<=x"0200000010";
mem(287)<=x"230000003a";
mem(288)<=x"0200000010";
mem(289)<=x"010000002f";
mem(290)<=x"5100000265";
mem(291)<=x"230000000a";
mem(292)<=x"0200000010";
mem(293)<=x"5200000000";
mem(294)<=x"2100000004";
mem(295)<=x"0200000029";
mem(296)<=x"2300000050";
mem(297)<=x"0200000010";
mem(298)<=x"2300000077";
mem(299)<=x"0200000010";
mem(300)<=x"230000006d";
mem(301)<=x"0200000010";
mem(302)<=x"2300000020";
mem(303)<=x"0200000010";
mem(304)<=x"230000004f";
mem(305)<=x"0200000010";
mem(306)<=x"2300000070";
mem(307)<=x"0200000010";
mem(308)<=x"2300000065";
mem(309)<=x"0200000010";
mem(310)<=x"230000006e";
mem(311)<=x"0200000010";
mem(312)<=x"230000003a";
mem(313)<=x"0200000010";
mem(314)<=x"2300000020";
mem(315)<=x"0200000010";
mem(316)<=x"010000002b";
mem(317)<=x"2200000005";
mem(318)<=x"230000000f";
mem(319)<=x"2200000006";
mem(320)<=x"2300000030";
mem(321)<=x"2200000007";
mem(322)<=x"2100000005";
mem(323)<=x"3800000000";
mem(324)<=x"3800000000";
mem(325)<=x"3800000000";
mem(326)<=x"3200000006";
mem(327)<=x"3100000007";
mem(328)<=x"0200000010";
mem(329)<=x"2100000005";
mem(330)<=x"3800000000";
mem(331)<=x"3800000000";
mem(332)<=x"3200000006";
mem(333)<=x"3100000007";
mem(334)<=x"0200000010";
mem(335)<=x"2100000005";
mem(336)<=x"3800000000";
mem(337)<=x"3200000006";
mem(338)<=x"3100000007";
mem(339)<=x"0200000010";
mem(340)<=x"2100000005";
mem(341)<=x"3200000006";
mem(342)<=x"3100000007";
mem(343)<=x"0200000010";
mem(344)<=x"2300000020";
mem(345)<=x"0200000010";
mem(346)<=x"010000002a";
mem(347)<=x"2200000005";
mem(348)<=x"2100000005";
mem(349)<=x"3800000000";
mem(350)<=x"3800000000";
mem(351)<=x"3800000000";
mem(352)<=x"3800000000";
mem(353)<=x"3800000000";
mem(354)<=x"3800000000";
mem(355)<=x"3800000000";
mem(356)<=x"3200000006";
mem(357)<=x"3100000007";
mem(358)<=x"0200000010";
mem(359)<=x"2100000005";
mem(360)<=x"3800000000";
mem(361)<=x"3800000000";
mem(362)<=x"3800000000";
mem(363)<=x"3800000000";
mem(364)<=x"3800000000";
mem(365)<=x"3800000000";
mem(366)<=x"3200000006";
mem(367)<=x"3100000007";
mem(368)<=x"0200000010";
mem(369)<=x"2100000005";
mem(370)<=x"3800000000";
mem(371)<=x"3800000000";
mem(372)<=x"3800000000";
mem(373)<=x"3800000000";
mem(374)<=x"3800000000";
mem(375)<=x"3200000006";
mem(376)<=x"3100000007";
mem(377)<=x"0200000010";
mem(378)<=x"2100000005";
mem(379)<=x"3800000000";
mem(380)<=x"3800000000";
mem(381)<=x"3800000000";
mem(382)<=x"3800000000";
mem(383)<=x"3200000006";
mem(384)<=x"3100000007";
mem(385)<=x"0200000010";
mem(386)<=x"2300000020";
mem(387)<=x"0200000010";
mem(388)<=x"2100000005";
mem(389)<=x"3800000000";
mem(390)<=x"3800000000";
mem(391)<=x"3800000000";
mem(392)<=x"3200000006";
mem(393)<=x"3100000007";
mem(394)<=x"0200000010";
mem(395)<=x"2100000005";
mem(396)<=x"3800000000";
mem(397)<=x"3800000000";
mem(398)<=x"3200000006";
mem(399)<=x"3100000007";
mem(400)<=x"0200000010";
mem(401)<=x"2100000005";
mem(402)<=x"3800000000";
mem(403)<=x"3200000006";
mem(404)<=x"3100000007";
mem(405)<=x"0200000010";
mem(406)<=x"2100000005";
mem(407)<=x"3200000006";
mem(408)<=x"3100000007";
mem(409)<=x"0200000010";
mem(410)<=x"230000000a";
mem(411)<=x"0200000010";
mem(412)<=x"5200000000";
mem(413)<=x"2300000050";
mem(414)<=x"0200000010";
mem(415)<=x"230000006c";
mem(416)<=x"0200000010";
mem(417)<=x"2300000065";
mem(418)<=x"0200000010";
mem(419)<=x"2300000061";
mem(420)<=x"0200000010";
mem(421)<=x"2300000073";
mem(422)<=x"0200000010";
mem(423)<=x"2300000065";
mem(424)<=x"0200000010";
mem(425)<=x"2300000020";
mem(426)<=x"0200000010";
mem(427)<=x"2300000049";
mem(428)<=x"0200000010";
mem(429)<=x"230000006e";
mem(430)<=x"0200000010";
mem(431)<=x"2300000070";
mem(432)<=x"0200000010";
mem(433)<=x"2300000075";
mem(434)<=x"0200000010";
mem(435)<=x"2300000074";
mem(436)<=x"0200000010";
mem(437)<=x"2300000020";
mem(438)<=x"0200000010";
mem(439)<=x"2300000063";
mem(440)<=x"0200000010";
mem(441)<=x"230000006d";
mem(442)<=x"0200000010";
mem(443)<=x"2300000064";
mem(444)<=x"0200000010";
mem(445)<=x"230000002e";
mem(446)<=x"0200000010";
mem(447)<=x"230000000a";
mem(448)<=x"0200000010";
mem(449)<=x"5200000000";
mem(450)<=x"010000002c";
mem(451)<=x"2200000005";
mem(452)<=x"13000001c6";
mem(453)<=x"5200000000";
mem(454)<=x"230000004d";
mem(455)<=x"0200000010";
mem(456)<=x"230000004f";
mem(457)<=x"0200000010";
mem(458)<=x"2300000053";
mem(459)<=x"0200000010";
mem(460)<=x"2300000020";
mem(461)<=x"0200000010";
mem(462)<=x"2300000045";
mem(463)<=x"0200000010";
mem(464)<=x"2300000052";
mem(465)<=x"0200000010";
mem(466)<=x"2300000052";
mem(467)<=x"0200000010";
mem(468)<=x"230000003a";
mem(469)<=x"0200000010";
mem(470)<=x"2300000001";
mem(471)<=x"2200000006";
mem(472)<=x"2300000030";
mem(473)<=x"2200000007";
mem(474)<=x"2100000005";
mem(475)<=x"3600000000";
mem(476)<=x"3600000000";
mem(477)<=x"3600000000";
mem(478)<=x"3600000000";
mem(479)<=x"3600000000";
mem(480)<=x"3200000006";
mem(481)<=x"3100000007";
mem(482)<=x"0200000010";
mem(483)<=x"2100000005";
mem(484)<=x"3600000000";
mem(485)<=x"3600000000";
mem(486)<=x"3600000000";
mem(487)<=x"3600000000";
mem(488)<=x"3200000006";
mem(489)<=x"3100000007";
mem(490)<=x"0200000010";
mem(491)<=x"2100000005";
mem(492)<=x"3600000000";
mem(493)<=x"3600000000";
mem(494)<=x"3600000000";
mem(495)<=x"3200000006";
mem(496)<=x"3100000007";
mem(497)<=x"0200000010";
mem(498)<=x"2100000005";
mem(499)<=x"3600000000";
mem(500)<=x"3600000000";
mem(501)<=x"3200000006";
mem(502)<=x"3100000007";
mem(503)<=x"0200000010";
mem(504)<=x"2100000005";
mem(505)<=x"3600000000";
mem(506)<=x"3200000006";
mem(507)<=x"3100000007";
mem(508)<=x"0200000010";
mem(509)<=x"2100000005";
mem(510)<=x"3200000006";
mem(511)<=x"3100000007";
mem(512)<=x"0200000010";
mem(513)<=x"230000000a";
mem(514)<=x"0200000010";
mem(515)<=x"5200000000";
mem(516)<=x"2300000054";
mem(517)<=x"0200000010";
mem(518)<=x"2300000031";
mem(519)<=x"0200000010";
mem(520)<=x"230000003a";
mem(521)<=x"0200000010";
mem(522)<=x"0100000024";
mem(523)<=x"5100000265";
mem(524)<=x"2300000075";
mem(525)<=x"0200000010";
mem(526)<=x"2300000073";
mem(527)<=x"0200000010";
mem(528)<=x"230000003b";
mem(529)<=x"0200000010";
mem(530)<=x"2300000054";
mem(531)<=x"0200000010";
mem(532)<=x"2300000032";
mem(533)<=x"0200000010";
mem(534)<=x"230000003a";
mem(535)<=x"0200000010";
mem(536)<=x"0100000025";
mem(537)<=x"5100000265";
mem(538)<=x"2300000075";
mem(539)<=x"0200000010";
mem(540)<=x"2300000073";
mem(541)<=x"0200000010";
mem(542)<=x"230000003b";
mem(543)<=x"0200000010";
mem(544)<=x"2300000054";
mem(545)<=x"0200000010";
mem(546)<=x"2300000033";
mem(547)<=x"0200000010";
mem(548)<=x"230000003a";
mem(549)<=x"0200000010";
mem(550)<=x"0100000026";
mem(551)<=x"5100000265";
mem(552)<=x"2300000075";
mem(553)<=x"0200000010";
mem(554)<=x"2300000073";
mem(555)<=x"0200000010";
mem(556)<=x"230000002e";
mem(557)<=x"0200000010";
mem(558)<=x"230000000a";
mem(559)<=x"0200000010";
mem(560)<=x"5200000000";
mem(561)<=x"2300000049";
mem(562)<=x"0200000010";
mem(563)<=x"2300000020";
mem(564)<=x"0200000010";
mem(565)<=x"2300000064";
mem(566)<=x"0200000010";
mem(567)<=x"230000006f";
mem(568)<=x"0200000010";
mem(569)<=x"230000006e";
mem(570)<=x"0200000010";
mem(571)<=x"2300000060";
mem(572)<=x"0200000010";
mem(573)<=x"2300000074";
mem(574)<=x"0200000010";
mem(575)<=x"2300000020";
mem(576)<=x"0200000010";
mem(577)<=x"230000006b";
mem(578)<=x"0200000010";
mem(579)<=x"230000006e";
mem(580)<=x"0200000010";
mem(581)<=x"230000006f";
mem(582)<=x"0200000010";
mem(583)<=x"2300000077";
mem(584)<=x"0200000010";
mem(585)<=x"2300000020";
mem(586)<=x"0200000010";
mem(587)<=x"2300000079";
mem(588)<=x"0200000010";
mem(589)<=x"230000006f";
mem(590)<=x"0200000010";
mem(591)<=x"2300000075";
mem(592)<=x"0200000010";
mem(593)<=x"2300000072";
mem(594)<=x"0200000010";
mem(595)<=x"2300000020";
mem(596)<=x"0200000010";
mem(597)<=x"2300000063";
mem(598)<=x"0200000010";
mem(599)<=x"230000006d";
mem(600)<=x"0200000010";
mem(601)<=x"2300000064";
mem(602)<=x"0200000010";
mem(603)<=x"230000000a";
mem(604)<=x"0200000010";
mem(605)<=x"5200000000";
mem(606)<=x"2300000010";
mem(607)<=x"2200000005";
mem(608)<=x"0100000013";
mem(609)<=x"3200000005";
mem(610)<=x"1300000260";
mem(611)<=x"0100000011";
mem(612)<=x"5200000000";
mem(613)<=x"0200000021";
mem(614)<=x"4100000020";
mem(615)<=x"0100000023";
mem(616)<=x"2200000005";
mem(617)<=x"230000000f";
mem(618)<=x"2200000006";
mem(619)<=x"2300000030";
mem(620)<=x"2200000007";
mem(621)<=x"2100000005";
mem(622)<=x"3800000000";
mem(623)<=x"3800000000";
mem(624)<=x"3800000000";
mem(625)<=x"3800000000";
mem(626)<=x"3200000006";
mem(627)<=x"3100000007";
mem(628)<=x"0200000010";
mem(629)<=x"2100000005";
mem(630)<=x"3800000000";
mem(631)<=x"3800000000";
mem(632)<=x"3800000000";
mem(633)<=x"3200000006";
mem(634)<=x"3100000007";
mem(635)<=x"0200000010";
mem(636)<=x"2100000005";
mem(637)<=x"3800000000";
mem(638)<=x"3800000000";
mem(639)<=x"3200000006";
mem(640)<=x"3100000007";
mem(641)<=x"0200000010";
mem(642)<=x"2100000005";
mem(643)<=x"3800000000";
mem(644)<=x"3200000006";
mem(645)<=x"3100000007";
mem(646)<=x"0200000010";
mem(647)<=x"2100000005";
mem(648)<=x"3200000006";
mem(649)<=x"3100000007";
mem(650)<=x"0200000010";
mem(651)<=x"5200000000";






end Behavioral;